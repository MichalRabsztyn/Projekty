1
0
48
6
54
27
31
18
50
64
7
33
62
